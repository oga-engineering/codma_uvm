// Simple declaration of the CPU VC sequencer.
typedef uvm_sequencer #(cpu_instruction) cpu_sequencer;