// TO be written: coverage file