typedef uvm_sequencer #(cpu_instruction) cpu_sequencer;