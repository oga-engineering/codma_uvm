package mem_pkg;

   `include "uvm_macros.svh"
   import uvm_pkg::*;

   `include "../uvcs/mem/mem_transaction.sv"
   `include "../uvcs/mem/mem_sequences.sv"
   `include "../uvcs/mem/mem_sequencer.sv"
   `include "../uvcs/mem/mem_driver.sv"
   `include "../uvcs/mem/mem_agent.sv"

endpackage